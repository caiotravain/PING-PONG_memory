// audio_nios.v

// Generated using ACDS version 16.1 196

`timescale 1 ps / 1 ps
module audio_nios (
		output wire        altpll_audio_locked_export,         //         altpll_audio_locked.export
		output wire        audio_conduit_end_XCK,              //           audio_conduit_end.XCK
		input  wire        audio_conduit_end_ADCDAT,           //                            .ADCDAT
		input  wire        audio_conduit_end_ADCLRC,           //                            .ADCLRC
		output wire        audio_conduit_end_DACDAT,           //                            .DACDAT
		input  wire        audio_conduit_end_DACLRC,           //                            .DACLRC
		input  wire        audio_conduit_end_BCLK,             //                            .BCLK
		input  wire        clk_clk,                            //                         clk.clk
		output wire        i2c_scl_external_connection_export, // i2c_scl_external_connection.export
		inout  wire        i2c_sda_external_connection_export, // i2c_sda_external_connection.export
		input  wire [3:0]  key_external_connection_export,     //     key_external_connection.export
		output wire [9:0]  pio_0_external_connection_export,   //   pio_0_external_connection.export
		output wire        pll_locked_export,                  //                  pll_locked.export
		output wire        pll_sdam_clk,                       //                    pll_sdam.clk
		input  wire        reset_reset_n,                      //                       reset.reset_n
		output wire [12:0] sdram_wire_addr,                    //                  sdram_wire.addr
		output wire [1:0]  sdram_wire_ba,                      //                            .ba
		output wire        sdram_wire_cas_n,                   //                            .cas_n
		output wire        sdram_wire_cke,                     //                            .cke
		output wire        sdram_wire_cs_n,                    //                            .cs_n
		inout  wire [15:0] sdram_wire_dq,                      //                            .dq
		output wire [1:0]  sdram_wire_dqm,                     //                            .dqm
		output wire        sdram_wire_ras_n,                   //                            .ras_n
		output wire        sdram_wire_we_n,                    //                            .we_n
		output wire [47:0] seg7_conduit_end_export,            //            seg7_conduit_end.export
		input  wire [9:0]  sw_external_connection_export       //      sw_external_connection.export
	);

	wire         pll_outclk0_clk;                                            // pll:outclk_0 -> [cpu_peripheral_bridge:s0_clk, irq_mapper:clk, irq_synchronizer:sender_clk, irq_synchronizer_001:sender_clk, jtag_uart:clk, mm_interconnect_0:pll_outclk0_clk, nios2_gen2_0:clk, onchip_memory2:clk, rst_controller_002:clk, rst_controller_003:clk, sdram:clk, sysid_qsys:clock, timer:clk]
	wire         altpll_audio_outclk0_clk;                                   // altpll_audio:outclk_0 -> [audio:avs_s1_clk, mm_interconnect_0:altpll_audio_outclk0_clk, rst_controller:clk]
	wire         pll_outclk2_clk;                                            // pll:outclk_2 -> [cpu_peripheral_bridge:m0_clk, i2c_scl:clk, i2c_sda:clk, irq_synchronizer:receiver_clk, irq_synchronizer_001:receiver_clk, key:clk, mm_interconnect_1:pll_outclk2_clk, pio_led:clk, rst_controller_001:clk, seg7:s_clk, sw:clk]
	wire  [31:0] nios2_gen2_0_data_master_readdata;                          // mm_interconnect_0:nios2_gen2_0_data_master_readdata -> nios2_gen2_0:d_readdata
	wire         nios2_gen2_0_data_master_waitrequest;                       // mm_interconnect_0:nios2_gen2_0_data_master_waitrequest -> nios2_gen2_0:d_waitrequest
	wire         nios2_gen2_0_data_master_debugaccess;                       // nios2_gen2_0:debug_mem_slave_debugaccess_to_roms -> mm_interconnect_0:nios2_gen2_0_data_master_debugaccess
	wire  [26:0] nios2_gen2_0_data_master_address;                           // nios2_gen2_0:d_address -> mm_interconnect_0:nios2_gen2_0_data_master_address
	wire   [3:0] nios2_gen2_0_data_master_byteenable;                        // nios2_gen2_0:d_byteenable -> mm_interconnect_0:nios2_gen2_0_data_master_byteenable
	wire         nios2_gen2_0_data_master_read;                              // nios2_gen2_0:d_read -> mm_interconnect_0:nios2_gen2_0_data_master_read
	wire         nios2_gen2_0_data_master_readdatavalid;                     // mm_interconnect_0:nios2_gen2_0_data_master_readdatavalid -> nios2_gen2_0:d_readdatavalid
	wire         nios2_gen2_0_data_master_write;                             // nios2_gen2_0:d_write -> mm_interconnect_0:nios2_gen2_0_data_master_write
	wire  [31:0] nios2_gen2_0_data_master_writedata;                         // nios2_gen2_0:d_writedata -> mm_interconnect_0:nios2_gen2_0_data_master_writedata
	wire  [31:0] nios2_gen2_0_instruction_master_readdata;                   // mm_interconnect_0:nios2_gen2_0_instruction_master_readdata -> nios2_gen2_0:i_readdata
	wire         nios2_gen2_0_instruction_master_waitrequest;                // mm_interconnect_0:nios2_gen2_0_instruction_master_waitrequest -> nios2_gen2_0:i_waitrequest
	wire  [26:0] nios2_gen2_0_instruction_master_address;                    // nios2_gen2_0:i_address -> mm_interconnect_0:nios2_gen2_0_instruction_master_address
	wire         nios2_gen2_0_instruction_master_read;                       // nios2_gen2_0:i_read -> mm_interconnect_0:nios2_gen2_0_instruction_master_read
	wire         nios2_gen2_0_instruction_master_readdatavalid;              // mm_interconnect_0:nios2_gen2_0_instruction_master_readdatavalid -> nios2_gen2_0:i_readdatavalid
	wire         mm_interconnect_0_jtag_uart_avalon_jtag_slave_chipselect;   // mm_interconnect_0:jtag_uart_avalon_jtag_slave_chipselect -> jtag_uart:av_chipselect
	wire  [31:0] mm_interconnect_0_jtag_uart_avalon_jtag_slave_readdata;     // jtag_uart:av_readdata -> mm_interconnect_0:jtag_uart_avalon_jtag_slave_readdata
	wire         mm_interconnect_0_jtag_uart_avalon_jtag_slave_waitrequest;  // jtag_uart:av_waitrequest -> mm_interconnect_0:jtag_uart_avalon_jtag_slave_waitrequest
	wire   [0:0] mm_interconnect_0_jtag_uart_avalon_jtag_slave_address;      // mm_interconnect_0:jtag_uart_avalon_jtag_slave_address -> jtag_uart:av_address
	wire         mm_interconnect_0_jtag_uart_avalon_jtag_slave_read;         // mm_interconnect_0:jtag_uart_avalon_jtag_slave_read -> jtag_uart:av_read_n
	wire         mm_interconnect_0_jtag_uart_avalon_jtag_slave_write;        // mm_interconnect_0:jtag_uart_avalon_jtag_slave_write -> jtag_uart:av_write_n
	wire  [31:0] mm_interconnect_0_jtag_uart_avalon_jtag_slave_writedata;    // mm_interconnect_0:jtag_uart_avalon_jtag_slave_writedata -> jtag_uart:av_writedata
	wire  [15:0] mm_interconnect_0_audio_avalon_slave_readdata;              // audio:avs_s1_readdata -> mm_interconnect_0:audio_avalon_slave_readdata
	wire   [2:0] mm_interconnect_0_audio_avalon_slave_address;               // mm_interconnect_0:audio_avalon_slave_address -> audio:avs_s1_address
	wire         mm_interconnect_0_audio_avalon_slave_read;                  // mm_interconnect_0:audio_avalon_slave_read -> audio:avs_s1_read
	wire         mm_interconnect_0_audio_avalon_slave_write;                 // mm_interconnect_0:audio_avalon_slave_write -> audio:avs_s1_write
	wire  [15:0] mm_interconnect_0_audio_avalon_slave_writedata;             // mm_interconnect_0:audio_avalon_slave_writedata -> audio:avs_s1_writedata
	wire  [31:0] mm_interconnect_0_sysid_qsys_control_slave_readdata;        // sysid_qsys:readdata -> mm_interconnect_0:sysid_qsys_control_slave_readdata
	wire   [0:0] mm_interconnect_0_sysid_qsys_control_slave_address;         // mm_interconnect_0:sysid_qsys_control_slave_address -> sysid_qsys:address
	wire  [31:0] mm_interconnect_0_nios2_gen2_0_debug_mem_slave_readdata;    // nios2_gen2_0:debug_mem_slave_readdata -> mm_interconnect_0:nios2_gen2_0_debug_mem_slave_readdata
	wire         mm_interconnect_0_nios2_gen2_0_debug_mem_slave_waitrequest; // nios2_gen2_0:debug_mem_slave_waitrequest -> mm_interconnect_0:nios2_gen2_0_debug_mem_slave_waitrequest
	wire         mm_interconnect_0_nios2_gen2_0_debug_mem_slave_debugaccess; // mm_interconnect_0:nios2_gen2_0_debug_mem_slave_debugaccess -> nios2_gen2_0:debug_mem_slave_debugaccess
	wire   [8:0] mm_interconnect_0_nios2_gen2_0_debug_mem_slave_address;     // mm_interconnect_0:nios2_gen2_0_debug_mem_slave_address -> nios2_gen2_0:debug_mem_slave_address
	wire         mm_interconnect_0_nios2_gen2_0_debug_mem_slave_read;        // mm_interconnect_0:nios2_gen2_0_debug_mem_slave_read -> nios2_gen2_0:debug_mem_slave_read
	wire   [3:0] mm_interconnect_0_nios2_gen2_0_debug_mem_slave_byteenable;  // mm_interconnect_0:nios2_gen2_0_debug_mem_slave_byteenable -> nios2_gen2_0:debug_mem_slave_byteenable
	wire         mm_interconnect_0_nios2_gen2_0_debug_mem_slave_write;       // mm_interconnect_0:nios2_gen2_0_debug_mem_slave_write -> nios2_gen2_0:debug_mem_slave_write
	wire  [31:0] mm_interconnect_0_nios2_gen2_0_debug_mem_slave_writedata;   // mm_interconnect_0:nios2_gen2_0_debug_mem_slave_writedata -> nios2_gen2_0:debug_mem_slave_writedata
	wire  [31:0] mm_interconnect_0_cpu_peripheral_bridge_s0_readdata;        // cpu_peripheral_bridge:s0_readdata -> mm_interconnect_0:cpu_peripheral_bridge_s0_readdata
	wire         mm_interconnect_0_cpu_peripheral_bridge_s0_waitrequest;     // cpu_peripheral_bridge:s0_waitrequest -> mm_interconnect_0:cpu_peripheral_bridge_s0_waitrequest
	wire         mm_interconnect_0_cpu_peripheral_bridge_s0_debugaccess;     // mm_interconnect_0:cpu_peripheral_bridge_s0_debugaccess -> cpu_peripheral_bridge:s0_debugaccess
	wire   [8:0] mm_interconnect_0_cpu_peripheral_bridge_s0_address;         // mm_interconnect_0:cpu_peripheral_bridge_s0_address -> cpu_peripheral_bridge:s0_address
	wire         mm_interconnect_0_cpu_peripheral_bridge_s0_read;            // mm_interconnect_0:cpu_peripheral_bridge_s0_read -> cpu_peripheral_bridge:s0_read
	wire   [3:0] mm_interconnect_0_cpu_peripheral_bridge_s0_byteenable;      // mm_interconnect_0:cpu_peripheral_bridge_s0_byteenable -> cpu_peripheral_bridge:s0_byteenable
	wire         mm_interconnect_0_cpu_peripheral_bridge_s0_readdatavalid;   // cpu_peripheral_bridge:s0_readdatavalid -> mm_interconnect_0:cpu_peripheral_bridge_s0_readdatavalid
	wire         mm_interconnect_0_cpu_peripheral_bridge_s0_write;           // mm_interconnect_0:cpu_peripheral_bridge_s0_write -> cpu_peripheral_bridge:s0_write
	wire  [31:0] mm_interconnect_0_cpu_peripheral_bridge_s0_writedata;       // mm_interconnect_0:cpu_peripheral_bridge_s0_writedata -> cpu_peripheral_bridge:s0_writedata
	wire   [0:0] mm_interconnect_0_cpu_peripheral_bridge_s0_burstcount;      // mm_interconnect_0:cpu_peripheral_bridge_s0_burstcount -> cpu_peripheral_bridge:s0_burstcount
	wire         mm_interconnect_0_onchip_memory2_s1_chipselect;             // mm_interconnect_0:onchip_memory2_s1_chipselect -> onchip_memory2:chipselect
	wire  [31:0] mm_interconnect_0_onchip_memory2_s1_readdata;               // onchip_memory2:readdata -> mm_interconnect_0:onchip_memory2_s1_readdata
	wire  [16:0] mm_interconnect_0_onchip_memory2_s1_address;                // mm_interconnect_0:onchip_memory2_s1_address -> onchip_memory2:address
	wire   [3:0] mm_interconnect_0_onchip_memory2_s1_byteenable;             // mm_interconnect_0:onchip_memory2_s1_byteenable -> onchip_memory2:byteenable
	wire         mm_interconnect_0_onchip_memory2_s1_write;                  // mm_interconnect_0:onchip_memory2_s1_write -> onchip_memory2:write
	wire  [31:0] mm_interconnect_0_onchip_memory2_s1_writedata;              // mm_interconnect_0:onchip_memory2_s1_writedata -> onchip_memory2:writedata
	wire         mm_interconnect_0_onchip_memory2_s1_clken;                  // mm_interconnect_0:onchip_memory2_s1_clken -> onchip_memory2:clken
	wire         mm_interconnect_0_timer_s1_chipselect;                      // mm_interconnect_0:timer_s1_chipselect -> timer:chipselect
	wire  [15:0] mm_interconnect_0_timer_s1_readdata;                        // timer:readdata -> mm_interconnect_0:timer_s1_readdata
	wire   [2:0] mm_interconnect_0_timer_s1_address;                         // mm_interconnect_0:timer_s1_address -> timer:address
	wire         mm_interconnect_0_timer_s1_write;                           // mm_interconnect_0:timer_s1_write -> timer:write_n
	wire  [15:0] mm_interconnect_0_timer_s1_writedata;                       // mm_interconnect_0:timer_s1_writedata -> timer:writedata
	wire         mm_interconnect_0_sdram_s1_chipselect;                      // mm_interconnect_0:sdram_s1_chipselect -> sdram:az_cs
	wire  [15:0] mm_interconnect_0_sdram_s1_readdata;                        // sdram:za_data -> mm_interconnect_0:sdram_s1_readdata
	wire         mm_interconnect_0_sdram_s1_waitrequest;                     // sdram:za_waitrequest -> mm_interconnect_0:sdram_s1_waitrequest
	wire  [24:0] mm_interconnect_0_sdram_s1_address;                         // mm_interconnect_0:sdram_s1_address -> sdram:az_addr
	wire         mm_interconnect_0_sdram_s1_read;                            // mm_interconnect_0:sdram_s1_read -> sdram:az_rd_n
	wire   [1:0] mm_interconnect_0_sdram_s1_byteenable;                      // mm_interconnect_0:sdram_s1_byteenable -> sdram:az_be_n
	wire         mm_interconnect_0_sdram_s1_readdatavalid;                   // sdram:za_valid -> mm_interconnect_0:sdram_s1_readdatavalid
	wire         mm_interconnect_0_sdram_s1_write;                           // mm_interconnect_0:sdram_s1_write -> sdram:az_wr_n
	wire  [15:0] mm_interconnect_0_sdram_s1_writedata;                       // mm_interconnect_0:sdram_s1_writedata -> sdram:az_data
	wire         cpu_peripheral_bridge_m0_waitrequest;                       // mm_interconnect_1:cpu_peripheral_bridge_m0_waitrequest -> cpu_peripheral_bridge:m0_waitrequest
	wire  [31:0] cpu_peripheral_bridge_m0_readdata;                          // mm_interconnect_1:cpu_peripheral_bridge_m0_readdata -> cpu_peripheral_bridge:m0_readdata
	wire         cpu_peripheral_bridge_m0_debugaccess;                       // cpu_peripheral_bridge:m0_debugaccess -> mm_interconnect_1:cpu_peripheral_bridge_m0_debugaccess
	wire   [8:0] cpu_peripheral_bridge_m0_address;                           // cpu_peripheral_bridge:m0_address -> mm_interconnect_1:cpu_peripheral_bridge_m0_address
	wire         cpu_peripheral_bridge_m0_read;                              // cpu_peripheral_bridge:m0_read -> mm_interconnect_1:cpu_peripheral_bridge_m0_read
	wire   [3:0] cpu_peripheral_bridge_m0_byteenable;                        // cpu_peripheral_bridge:m0_byteenable -> mm_interconnect_1:cpu_peripheral_bridge_m0_byteenable
	wire         cpu_peripheral_bridge_m0_readdatavalid;                     // mm_interconnect_1:cpu_peripheral_bridge_m0_readdatavalid -> cpu_peripheral_bridge:m0_readdatavalid
	wire  [31:0] cpu_peripheral_bridge_m0_writedata;                         // cpu_peripheral_bridge:m0_writedata -> mm_interconnect_1:cpu_peripheral_bridge_m0_writedata
	wire         cpu_peripheral_bridge_m0_write;                             // cpu_peripheral_bridge:m0_write -> mm_interconnect_1:cpu_peripheral_bridge_m0_write
	wire   [0:0] cpu_peripheral_bridge_m0_burstcount;                        // cpu_peripheral_bridge:m0_burstcount -> mm_interconnect_1:cpu_peripheral_bridge_m0_burstcount
	wire   [7:0] mm_interconnect_1_seg7_avalon_slave_readdata;               // seg7:s_readdata -> mm_interconnect_1:seg7_avalon_slave_readdata
	wire   [2:0] mm_interconnect_1_seg7_avalon_slave_address;                // mm_interconnect_1:seg7_avalon_slave_address -> seg7:s_address
	wire         mm_interconnect_1_seg7_avalon_slave_read;                   // mm_interconnect_1:seg7_avalon_slave_read -> seg7:s_read
	wire         mm_interconnect_1_seg7_avalon_slave_write;                  // mm_interconnect_1:seg7_avalon_slave_write -> seg7:s_write
	wire   [7:0] mm_interconnect_1_seg7_avalon_slave_writedata;              // mm_interconnect_1:seg7_avalon_slave_writedata -> seg7:s_writedata
	wire         mm_interconnect_1_key_s1_chipselect;                        // mm_interconnect_1:key_s1_chipselect -> key:chipselect
	wire  [31:0] mm_interconnect_1_key_s1_readdata;                          // key:readdata -> mm_interconnect_1:key_s1_readdata
	wire   [1:0] mm_interconnect_1_key_s1_address;                           // mm_interconnect_1:key_s1_address -> key:address
	wire         mm_interconnect_1_key_s1_write;                             // mm_interconnect_1:key_s1_write -> key:write_n
	wire  [31:0] mm_interconnect_1_key_s1_writedata;                         // mm_interconnect_1:key_s1_writedata -> key:writedata
	wire         mm_interconnect_1_pio_led_s1_chipselect;                    // mm_interconnect_1:pio_led_s1_chipselect -> pio_led:chipselect
	wire  [31:0] mm_interconnect_1_pio_led_s1_readdata;                      // pio_led:readdata -> mm_interconnect_1:pio_led_s1_readdata
	wire   [1:0] mm_interconnect_1_pio_led_s1_address;                       // mm_interconnect_1:pio_led_s1_address -> pio_led:address
	wire         mm_interconnect_1_pio_led_s1_write;                         // mm_interconnect_1:pio_led_s1_write -> pio_led:write_n
	wire  [31:0] mm_interconnect_1_pio_led_s1_writedata;                     // mm_interconnect_1:pio_led_s1_writedata -> pio_led:writedata
	wire         mm_interconnect_1_sw_s1_chipselect;                         // mm_interconnect_1:sw_s1_chipselect -> sw:chipselect
	wire  [31:0] mm_interconnect_1_sw_s1_readdata;                           // sw:readdata -> mm_interconnect_1:sw_s1_readdata
	wire   [1:0] mm_interconnect_1_sw_s1_address;                            // mm_interconnect_1:sw_s1_address -> sw:address
	wire         mm_interconnect_1_sw_s1_write;                              // mm_interconnect_1:sw_s1_write -> sw:write_n
	wire  [31:0] mm_interconnect_1_sw_s1_writedata;                          // mm_interconnect_1:sw_s1_writedata -> sw:writedata
	wire         mm_interconnect_1_i2c_scl_s1_chipselect;                    // mm_interconnect_1:i2c_scl_s1_chipselect -> i2c_scl:chipselect
	wire  [31:0] mm_interconnect_1_i2c_scl_s1_readdata;                      // i2c_scl:readdata -> mm_interconnect_1:i2c_scl_s1_readdata
	wire   [1:0] mm_interconnect_1_i2c_scl_s1_address;                       // mm_interconnect_1:i2c_scl_s1_address -> i2c_scl:address
	wire         mm_interconnect_1_i2c_scl_s1_write;                         // mm_interconnect_1:i2c_scl_s1_write -> i2c_scl:write_n
	wire  [31:0] mm_interconnect_1_i2c_scl_s1_writedata;                     // mm_interconnect_1:i2c_scl_s1_writedata -> i2c_scl:writedata
	wire         mm_interconnect_1_i2c_sda_s1_chipselect;                    // mm_interconnect_1:i2c_sda_s1_chipselect -> i2c_sda:chipselect
	wire  [31:0] mm_interconnect_1_i2c_sda_s1_readdata;                      // i2c_sda:readdata -> mm_interconnect_1:i2c_sda_s1_readdata
	wire   [1:0] mm_interconnect_1_i2c_sda_s1_address;                       // mm_interconnect_1:i2c_sda_s1_address -> i2c_sda:address
	wire         mm_interconnect_1_i2c_sda_s1_write;                         // mm_interconnect_1:i2c_sda_s1_write -> i2c_sda:write_n
	wire  [31:0] mm_interconnect_1_i2c_sda_s1_writedata;                     // mm_interconnect_1:i2c_sda_s1_writedata -> i2c_sda:writedata
	wire         irq_mapper_receiver0_irq;                                   // timer:irq -> irq_mapper:receiver0_irq
	wire         irq_mapper_receiver1_irq;                                   // jtag_uart:av_irq -> irq_mapper:receiver1_irq
	wire  [31:0] nios2_gen2_0_irq_irq;                                       // irq_mapper:sender_irq -> nios2_gen2_0:irq
	wire         irq_mapper_receiver2_irq;                                   // irq_synchronizer:sender_irq -> irq_mapper:receiver2_irq
	wire   [0:0] irq_synchronizer_receiver_irq;                              // key:irq -> irq_synchronizer:receiver_irq
	wire         irq_mapper_receiver3_irq;                                   // irq_synchronizer_001:sender_irq -> irq_mapper:receiver3_irq
	wire   [0:0] irq_synchronizer_001_receiver_irq;                          // sw:irq -> irq_synchronizer_001:receiver_irq
	wire         rst_controller_reset_out_reset;                             // rst_controller:reset_out -> [audio:avs_s1_reset, mm_interconnect_0:audio_clock_sink_reset_reset_bridge_in_reset_reset]
	wire         rst_controller_001_reset_out_reset;                         // rst_controller_001:reset_out -> [cpu_peripheral_bridge:m0_reset, i2c_scl:reset_n, i2c_sda:reset_n, irq_synchronizer:receiver_reset, irq_synchronizer_001:receiver_reset, key:reset_n, mm_interconnect_1:cpu_peripheral_bridge_m0_reset_reset_bridge_in_reset_reset, pio_led:reset_n, seg7:s_reset, sw:reset_n]
	wire         rst_controller_002_reset_out_reset;                         // rst_controller_002:reset_out -> [cpu_peripheral_bridge:s0_reset, jtag_uart:rst_n, mm_interconnect_0:jtag_uart_reset_reset_bridge_in_reset_reset, onchip_memory2:reset, rst_translator:in_reset, sdram:reset_n, sysid_qsys:reset_n, timer:reset_n]
	wire         rst_controller_002_reset_out_reset_req;                     // rst_controller_002:reset_req -> [onchip_memory2:reset_req, rst_translator:reset_req_in]
	wire         rst_controller_003_reset_out_reset;                         // rst_controller_003:reset_out -> [irq_mapper:reset, irq_synchronizer:sender_reset, irq_synchronizer_001:sender_reset, mm_interconnect_0:nios2_gen2_0_reset_reset_bridge_in_reset_reset, nios2_gen2_0:reset_n, rst_translator_001:in_reset]
	wire         rst_controller_003_reset_out_reset_req;                     // rst_controller_003:reset_req -> [nios2_gen2_0:reset_req, rst_translator_001:reset_req_in]
	wire         nios2_gen2_0_debug_reset_request_reset;                     // nios2_gen2_0:debug_reset_request -> rst_controller_003:reset_in1

	audio_nios_altpll_audio altpll_audio (
		.refclk   (clk_clk),                    //  refclk.clk
		.rst      (~reset_reset_n),             //   reset.reset
		.outclk_0 (altpll_audio_outclk0_clk),   // outclk0.clk
		.locked   (altpll_audio_locked_export)  //  locked.export
	);

	AUDIO_IF audio (
		.avs_s1_address       (mm_interconnect_0_audio_avalon_slave_address),   //     avalon_slave.address
		.avs_s1_read          (mm_interconnect_0_audio_avalon_slave_read),      //                 .read
		.avs_s1_readdata      (mm_interconnect_0_audio_avalon_slave_readdata),  //                 .readdata
		.avs_s1_write         (mm_interconnect_0_audio_avalon_slave_write),     //                 .write
		.avs_s1_writedata     (mm_interconnect_0_audio_avalon_slave_writedata), //                 .writedata
		.avs_s1_clk           (altpll_audio_outclk0_clk),                       //       clock_sink.clk
		.avs_s1_reset         (rst_controller_reset_out_reset),                 // clock_sink_reset.reset
		.avs_s1_export_XCK    (audio_conduit_end_XCK),                          //      conduit_end.export
		.avs_s1_export_ADCDAT (audio_conduit_end_ADCDAT),                       //                 .export
		.avs_s1_export_ADCLRC (audio_conduit_end_ADCLRC),                       //                 .export
		.avs_s1_export_DACDAT (audio_conduit_end_DACDAT),                       //                 .export
		.avs_s1_export_DACLRC (audio_conduit_end_DACLRC),                       //                 .export
		.avs_s1_export_BCLK   (audio_conduit_end_BCLK)                          //                 .export
	);

	altera_avalon_mm_clock_crossing_bridge #(
		.DATA_WIDTH          (32),
		.SYMBOL_WIDTH        (8),
		.HDL_ADDR_WIDTH      (9),
		.BURSTCOUNT_WIDTH    (1),
		.COMMAND_FIFO_DEPTH  (32),
		.RESPONSE_FIFO_DEPTH (64),
		.MASTER_SYNC_DEPTH   (3),
		.SLAVE_SYNC_DEPTH    (3)
	) cpu_peripheral_bridge (
		.m0_clk           (pll_outclk2_clk),                                          //   m0_clk.clk
		.m0_reset         (rst_controller_001_reset_out_reset),                       // m0_reset.reset
		.s0_clk           (pll_outclk0_clk),                                          //   s0_clk.clk
		.s0_reset         (rst_controller_002_reset_out_reset),                       // s0_reset.reset
		.s0_waitrequest   (mm_interconnect_0_cpu_peripheral_bridge_s0_waitrequest),   //       s0.waitrequest
		.s0_readdata      (mm_interconnect_0_cpu_peripheral_bridge_s0_readdata),      //         .readdata
		.s0_readdatavalid (mm_interconnect_0_cpu_peripheral_bridge_s0_readdatavalid), //         .readdatavalid
		.s0_burstcount    (mm_interconnect_0_cpu_peripheral_bridge_s0_burstcount),    //         .burstcount
		.s0_writedata     (mm_interconnect_0_cpu_peripheral_bridge_s0_writedata),     //         .writedata
		.s0_address       (mm_interconnect_0_cpu_peripheral_bridge_s0_address),       //         .address
		.s0_write         (mm_interconnect_0_cpu_peripheral_bridge_s0_write),         //         .write
		.s0_read          (mm_interconnect_0_cpu_peripheral_bridge_s0_read),          //         .read
		.s0_byteenable    (mm_interconnect_0_cpu_peripheral_bridge_s0_byteenable),    //         .byteenable
		.s0_debugaccess   (mm_interconnect_0_cpu_peripheral_bridge_s0_debugaccess),   //         .debugaccess
		.m0_waitrequest   (cpu_peripheral_bridge_m0_waitrequest),                     //       m0.waitrequest
		.m0_readdata      (cpu_peripheral_bridge_m0_readdata),                        //         .readdata
		.m0_readdatavalid (cpu_peripheral_bridge_m0_readdatavalid),                   //         .readdatavalid
		.m0_burstcount    (cpu_peripheral_bridge_m0_burstcount),                      //         .burstcount
		.m0_writedata     (cpu_peripheral_bridge_m0_writedata),                       //         .writedata
		.m0_address       (cpu_peripheral_bridge_m0_address),                         //         .address
		.m0_write         (cpu_peripheral_bridge_m0_write),                           //         .write
		.m0_read          (cpu_peripheral_bridge_m0_read),                            //         .read
		.m0_byteenable    (cpu_peripheral_bridge_m0_byteenable),                      //         .byteenable
		.m0_debugaccess   (cpu_peripheral_bridge_m0_debugaccess)                      //         .debugaccess
	);

	audio_nios_i2c_scl i2c_scl (
		.clk        (pll_outclk2_clk),                         //                 clk.clk
		.reset_n    (~rst_controller_001_reset_out_reset),     //               reset.reset_n
		.address    (mm_interconnect_1_i2c_scl_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_1_i2c_scl_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_1_i2c_scl_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_1_i2c_scl_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_1_i2c_scl_s1_readdata),   //                    .readdata
		.out_port   (i2c_scl_external_connection_export)       // external_connection.export
	);

	audio_nios_i2c_sda i2c_sda (
		.clk        (pll_outclk2_clk),                         //                 clk.clk
		.reset_n    (~rst_controller_001_reset_out_reset),     //               reset.reset_n
		.address    (mm_interconnect_1_i2c_sda_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_1_i2c_sda_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_1_i2c_sda_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_1_i2c_sda_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_1_i2c_sda_s1_readdata),   //                    .readdata
		.bidir_port (i2c_sda_external_connection_export)       // external_connection.export
	);

	audio_nios_jtag_uart jtag_uart (
		.clk            (pll_outclk0_clk),                                           //               clk.clk
		.rst_n          (~rst_controller_002_reset_out_reset),                       //             reset.reset_n
		.av_chipselect  (mm_interconnect_0_jtag_uart_avalon_jtag_slave_chipselect),  // avalon_jtag_slave.chipselect
		.av_address     (mm_interconnect_0_jtag_uart_avalon_jtag_slave_address),     //                  .address
		.av_read_n      (~mm_interconnect_0_jtag_uart_avalon_jtag_slave_read),       //                  .read_n
		.av_readdata    (mm_interconnect_0_jtag_uart_avalon_jtag_slave_readdata),    //                  .readdata
		.av_write_n     (~mm_interconnect_0_jtag_uart_avalon_jtag_slave_write),      //                  .write_n
		.av_writedata   (mm_interconnect_0_jtag_uart_avalon_jtag_slave_writedata),   //                  .writedata
		.av_waitrequest (mm_interconnect_0_jtag_uart_avalon_jtag_slave_waitrequest), //                  .waitrequest
		.av_irq         (irq_mapper_receiver1_irq)                                   //               irq.irq
	);

	audio_nios_key key (
		.clk        (pll_outclk2_clk),                     //                 clk.clk
		.reset_n    (~rst_controller_001_reset_out_reset), //               reset.reset_n
		.address    (mm_interconnect_1_key_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_1_key_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_1_key_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_1_key_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_1_key_s1_readdata),   //                    .readdata
		.in_port    (key_external_connection_export),      // external_connection.export
		.irq        (irq_synchronizer_receiver_irq)        //                 irq.irq
	);

	audio_nios_nios2_gen2_0 nios2_gen2_0 (
		.clk                                 (pll_outclk0_clk),                                            //                       clk.clk
		.reset_n                             (~rst_controller_003_reset_out_reset),                        //                     reset.reset_n
		.reset_req                           (rst_controller_003_reset_out_reset_req),                     //                          .reset_req
		.d_address                           (nios2_gen2_0_data_master_address),                           //               data_master.address
		.d_byteenable                        (nios2_gen2_0_data_master_byteenable),                        //                          .byteenable
		.d_read                              (nios2_gen2_0_data_master_read),                              //                          .read
		.d_readdata                          (nios2_gen2_0_data_master_readdata),                          //                          .readdata
		.d_waitrequest                       (nios2_gen2_0_data_master_waitrequest),                       //                          .waitrequest
		.d_write                             (nios2_gen2_0_data_master_write),                             //                          .write
		.d_writedata                         (nios2_gen2_0_data_master_writedata),                         //                          .writedata
		.d_readdatavalid                     (nios2_gen2_0_data_master_readdatavalid),                     //                          .readdatavalid
		.debug_mem_slave_debugaccess_to_roms (nios2_gen2_0_data_master_debugaccess),                       //                          .debugaccess
		.i_address                           (nios2_gen2_0_instruction_master_address),                    //        instruction_master.address
		.i_read                              (nios2_gen2_0_instruction_master_read),                       //                          .read
		.i_readdata                          (nios2_gen2_0_instruction_master_readdata),                   //                          .readdata
		.i_waitrequest                       (nios2_gen2_0_instruction_master_waitrequest),                //                          .waitrequest
		.i_readdatavalid                     (nios2_gen2_0_instruction_master_readdatavalid),              //                          .readdatavalid
		.irq                                 (nios2_gen2_0_irq_irq),                                       //                       irq.irq
		.debug_reset_request                 (nios2_gen2_0_debug_reset_request_reset),                     //       debug_reset_request.reset
		.debug_mem_slave_address             (mm_interconnect_0_nios2_gen2_0_debug_mem_slave_address),     //           debug_mem_slave.address
		.debug_mem_slave_byteenable          (mm_interconnect_0_nios2_gen2_0_debug_mem_slave_byteenable),  //                          .byteenable
		.debug_mem_slave_debugaccess         (mm_interconnect_0_nios2_gen2_0_debug_mem_slave_debugaccess), //                          .debugaccess
		.debug_mem_slave_read                (mm_interconnect_0_nios2_gen2_0_debug_mem_slave_read),        //                          .read
		.debug_mem_slave_readdata            (mm_interconnect_0_nios2_gen2_0_debug_mem_slave_readdata),    //                          .readdata
		.debug_mem_slave_waitrequest         (mm_interconnect_0_nios2_gen2_0_debug_mem_slave_waitrequest), //                          .waitrequest
		.debug_mem_slave_write               (mm_interconnect_0_nios2_gen2_0_debug_mem_slave_write),       //                          .write
		.debug_mem_slave_writedata           (mm_interconnect_0_nios2_gen2_0_debug_mem_slave_writedata),   //                          .writedata
		.dummy_ci_port                       ()                                                            // custom_instruction_master.readra
	);

	audio_nios_onchip_memory2 onchip_memory2 (
		.clk        (pll_outclk0_clk),                                //   clk1.clk
		.address    (mm_interconnect_0_onchip_memory2_s1_address),    //     s1.address
		.clken      (mm_interconnect_0_onchip_memory2_s1_clken),      //       .clken
		.chipselect (mm_interconnect_0_onchip_memory2_s1_chipselect), //       .chipselect
		.write      (mm_interconnect_0_onchip_memory2_s1_write),      //       .write
		.readdata   (mm_interconnect_0_onchip_memory2_s1_readdata),   //       .readdata
		.writedata  (mm_interconnect_0_onchip_memory2_s1_writedata),  //       .writedata
		.byteenable (mm_interconnect_0_onchip_memory2_s1_byteenable), //       .byteenable
		.reset      (rst_controller_002_reset_out_reset),             // reset1.reset
		.reset_req  (rst_controller_002_reset_out_reset_req),         //       .reset_req
		.freeze     (1'b0)                                            // (terminated)
	);

	audio_nios_pio_led pio_led (
		.clk        (pll_outclk2_clk),                         //                 clk.clk
		.reset_n    (~rst_controller_001_reset_out_reset),     //               reset.reset_n
		.address    (mm_interconnect_1_pio_led_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_1_pio_led_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_1_pio_led_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_1_pio_led_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_1_pio_led_s1_readdata),   //                    .readdata
		.out_port   (pio_0_external_connection_export)         // external_connection.export
	);

	audio_nios_pll pll (
		.refclk   (clk_clk),           //  refclk.clk
		.rst      (~reset_reset_n),    //   reset.reset
		.outclk_0 (pll_outclk0_clk),   // outclk0.clk
		.outclk_1 (pll_sdam_clk),      // outclk1.clk
		.outclk_2 (pll_outclk2_clk),   // outclk2.clk
		.locked   (pll_locked_export)  //  locked.export
	);

	audio_nios_sdram sdram (
		.clk            (pll_outclk0_clk),                          //   clk.clk
		.reset_n        (~rst_controller_002_reset_out_reset),      // reset.reset_n
		.az_addr        (mm_interconnect_0_sdram_s1_address),       //    s1.address
		.az_be_n        (~mm_interconnect_0_sdram_s1_byteenable),   //      .byteenable_n
		.az_cs          (mm_interconnect_0_sdram_s1_chipselect),    //      .chipselect
		.az_data        (mm_interconnect_0_sdram_s1_writedata),     //      .writedata
		.az_rd_n        (~mm_interconnect_0_sdram_s1_read),         //      .read_n
		.az_wr_n        (~mm_interconnect_0_sdram_s1_write),        //      .write_n
		.za_data        (mm_interconnect_0_sdram_s1_readdata),      //      .readdata
		.za_valid       (mm_interconnect_0_sdram_s1_readdatavalid), //      .readdatavalid
		.za_waitrequest (mm_interconnect_0_sdram_s1_waitrequest),   //      .waitrequest
		.zs_addr        (sdram_wire_addr),                          //  wire.export
		.zs_ba          (sdram_wire_ba),                            //      .export
		.zs_cas_n       (sdram_wire_cas_n),                         //      .export
		.zs_cke         (sdram_wire_cke),                           //      .export
		.zs_cs_n        (sdram_wire_cs_n),                          //      .export
		.zs_dq          (sdram_wire_dq),                            //      .export
		.zs_dqm         (sdram_wire_dqm),                           //      .export
		.zs_ras_n       (sdram_wire_ras_n),                         //      .export
		.zs_we_n        (sdram_wire_we_n)                           //      .export
	);

	SEG7_IF #(
		.SEG7_NUM       (6),
		.ADDR_WIDTH     (3),
		.DEFAULT_ACTIVE (1),
		.LOW_ACTIVE     (1)
	) seg7 (
		.s_address   (mm_interconnect_1_seg7_avalon_slave_address),   //     avalon_slave.address
		.s_read      (mm_interconnect_1_seg7_avalon_slave_read),      //                 .read
		.s_readdata  (mm_interconnect_1_seg7_avalon_slave_readdata),  //                 .readdata
		.s_write     (mm_interconnect_1_seg7_avalon_slave_write),     //                 .write
		.s_writedata (mm_interconnect_1_seg7_avalon_slave_writedata), //                 .writedata
		.SEG7        (seg7_conduit_end_export),                       //      conduit_end.export
		.s_clk       (pll_outclk2_clk),                               //       clock_sink.clk
		.s_reset     (rst_controller_001_reset_out_reset)             // clock_sink_reset.reset
	);

	audio_nios_sw sw (
		.clk        (pll_outclk2_clk),                     //                 clk.clk
		.reset_n    (~rst_controller_001_reset_out_reset), //               reset.reset_n
		.address    (mm_interconnect_1_sw_s1_address),     //                  s1.address
		.write_n    (~mm_interconnect_1_sw_s1_write),      //                    .write_n
		.writedata  (mm_interconnect_1_sw_s1_writedata),   //                    .writedata
		.chipselect (mm_interconnect_1_sw_s1_chipselect),  //                    .chipselect
		.readdata   (mm_interconnect_1_sw_s1_readdata),    //                    .readdata
		.in_port    (sw_external_connection_export),       // external_connection.export
		.irq        (irq_synchronizer_001_receiver_irq)    //                 irq.irq
	);

	audio_nios_sysid_qsys sysid_qsys (
		.clock    (pll_outclk0_clk),                                     //           clk.clk
		.reset_n  (~rst_controller_002_reset_out_reset),                 //         reset.reset_n
		.readdata (mm_interconnect_0_sysid_qsys_control_slave_readdata), // control_slave.readdata
		.address  (mm_interconnect_0_sysid_qsys_control_slave_address)   //              .address
	);

	audio_nios_timer timer (
		.clk        (pll_outclk0_clk),                       //   clk.clk
		.reset_n    (~rst_controller_002_reset_out_reset),   // reset.reset_n
		.address    (mm_interconnect_0_timer_s1_address),    //    s1.address
		.writedata  (mm_interconnect_0_timer_s1_writedata),  //      .writedata
		.readdata   (mm_interconnect_0_timer_s1_readdata),   //      .readdata
		.chipselect (mm_interconnect_0_timer_s1_chipselect), //      .chipselect
		.write_n    (~mm_interconnect_0_timer_s1_write),     //      .write_n
		.irq        (irq_mapper_receiver0_irq)               //   irq.irq
	);

	audio_nios_mm_interconnect_0 mm_interconnect_0 (
		.altpll_audio_outclk0_clk                           (altpll_audio_outclk0_clk),                                   //                         altpll_audio_outclk0.clk
		.pll_outclk0_clk                                    (pll_outclk0_clk),                                            //                                  pll_outclk0.clk
		.audio_clock_sink_reset_reset_bridge_in_reset_reset (rst_controller_reset_out_reset),                             // audio_clock_sink_reset_reset_bridge_in_reset.reset
		.jtag_uart_reset_reset_bridge_in_reset_reset        (rst_controller_002_reset_out_reset),                         //        jtag_uart_reset_reset_bridge_in_reset.reset
		.nios2_gen2_0_reset_reset_bridge_in_reset_reset     (rst_controller_003_reset_out_reset),                         //     nios2_gen2_0_reset_reset_bridge_in_reset.reset
		.nios2_gen2_0_data_master_address                   (nios2_gen2_0_data_master_address),                           //                     nios2_gen2_0_data_master.address
		.nios2_gen2_0_data_master_waitrequest               (nios2_gen2_0_data_master_waitrequest),                       //                                             .waitrequest
		.nios2_gen2_0_data_master_byteenable                (nios2_gen2_0_data_master_byteenable),                        //                                             .byteenable
		.nios2_gen2_0_data_master_read                      (nios2_gen2_0_data_master_read),                              //                                             .read
		.nios2_gen2_0_data_master_readdata                  (nios2_gen2_0_data_master_readdata),                          //                                             .readdata
		.nios2_gen2_0_data_master_readdatavalid             (nios2_gen2_0_data_master_readdatavalid),                     //                                             .readdatavalid
		.nios2_gen2_0_data_master_write                     (nios2_gen2_0_data_master_write),                             //                                             .write
		.nios2_gen2_0_data_master_writedata                 (nios2_gen2_0_data_master_writedata),                         //                                             .writedata
		.nios2_gen2_0_data_master_debugaccess               (nios2_gen2_0_data_master_debugaccess),                       //                                             .debugaccess
		.nios2_gen2_0_instruction_master_address            (nios2_gen2_0_instruction_master_address),                    //              nios2_gen2_0_instruction_master.address
		.nios2_gen2_0_instruction_master_waitrequest        (nios2_gen2_0_instruction_master_waitrequest),                //                                             .waitrequest
		.nios2_gen2_0_instruction_master_read               (nios2_gen2_0_instruction_master_read),                       //                                             .read
		.nios2_gen2_0_instruction_master_readdata           (nios2_gen2_0_instruction_master_readdata),                   //                                             .readdata
		.nios2_gen2_0_instruction_master_readdatavalid      (nios2_gen2_0_instruction_master_readdatavalid),              //                                             .readdatavalid
		.audio_avalon_slave_address                         (mm_interconnect_0_audio_avalon_slave_address),               //                           audio_avalon_slave.address
		.audio_avalon_slave_write                           (mm_interconnect_0_audio_avalon_slave_write),                 //                                             .write
		.audio_avalon_slave_read                            (mm_interconnect_0_audio_avalon_slave_read),                  //                                             .read
		.audio_avalon_slave_readdata                        (mm_interconnect_0_audio_avalon_slave_readdata),              //                                             .readdata
		.audio_avalon_slave_writedata                       (mm_interconnect_0_audio_avalon_slave_writedata),             //                                             .writedata
		.cpu_peripheral_bridge_s0_address                   (mm_interconnect_0_cpu_peripheral_bridge_s0_address),         //                     cpu_peripheral_bridge_s0.address
		.cpu_peripheral_bridge_s0_write                     (mm_interconnect_0_cpu_peripheral_bridge_s0_write),           //                                             .write
		.cpu_peripheral_bridge_s0_read                      (mm_interconnect_0_cpu_peripheral_bridge_s0_read),            //                                             .read
		.cpu_peripheral_bridge_s0_readdata                  (mm_interconnect_0_cpu_peripheral_bridge_s0_readdata),        //                                             .readdata
		.cpu_peripheral_bridge_s0_writedata                 (mm_interconnect_0_cpu_peripheral_bridge_s0_writedata),       //                                             .writedata
		.cpu_peripheral_bridge_s0_burstcount                (mm_interconnect_0_cpu_peripheral_bridge_s0_burstcount),      //                                             .burstcount
		.cpu_peripheral_bridge_s0_byteenable                (mm_interconnect_0_cpu_peripheral_bridge_s0_byteenable),      //                                             .byteenable
		.cpu_peripheral_bridge_s0_readdatavalid             (mm_interconnect_0_cpu_peripheral_bridge_s0_readdatavalid),   //                                             .readdatavalid
		.cpu_peripheral_bridge_s0_waitrequest               (mm_interconnect_0_cpu_peripheral_bridge_s0_waitrequest),     //                                             .waitrequest
		.cpu_peripheral_bridge_s0_debugaccess               (mm_interconnect_0_cpu_peripheral_bridge_s0_debugaccess),     //                                             .debugaccess
		.jtag_uart_avalon_jtag_slave_address                (mm_interconnect_0_jtag_uart_avalon_jtag_slave_address),      //                  jtag_uart_avalon_jtag_slave.address
		.jtag_uart_avalon_jtag_slave_write                  (mm_interconnect_0_jtag_uart_avalon_jtag_slave_write),        //                                             .write
		.jtag_uart_avalon_jtag_slave_read                   (mm_interconnect_0_jtag_uart_avalon_jtag_slave_read),         //                                             .read
		.jtag_uart_avalon_jtag_slave_readdata               (mm_interconnect_0_jtag_uart_avalon_jtag_slave_readdata),     //                                             .readdata
		.jtag_uart_avalon_jtag_slave_writedata              (mm_interconnect_0_jtag_uart_avalon_jtag_slave_writedata),    //                                             .writedata
		.jtag_uart_avalon_jtag_slave_waitrequest            (mm_interconnect_0_jtag_uart_avalon_jtag_slave_waitrequest),  //                                             .waitrequest
		.jtag_uart_avalon_jtag_slave_chipselect             (mm_interconnect_0_jtag_uart_avalon_jtag_slave_chipselect),   //                                             .chipselect
		.nios2_gen2_0_debug_mem_slave_address               (mm_interconnect_0_nios2_gen2_0_debug_mem_slave_address),     //                 nios2_gen2_0_debug_mem_slave.address
		.nios2_gen2_0_debug_mem_slave_write                 (mm_interconnect_0_nios2_gen2_0_debug_mem_slave_write),       //                                             .write
		.nios2_gen2_0_debug_mem_slave_read                  (mm_interconnect_0_nios2_gen2_0_debug_mem_slave_read),        //                                             .read
		.nios2_gen2_0_debug_mem_slave_readdata              (mm_interconnect_0_nios2_gen2_0_debug_mem_slave_readdata),    //                                             .readdata
		.nios2_gen2_0_debug_mem_slave_writedata             (mm_interconnect_0_nios2_gen2_0_debug_mem_slave_writedata),   //                                             .writedata
		.nios2_gen2_0_debug_mem_slave_byteenable            (mm_interconnect_0_nios2_gen2_0_debug_mem_slave_byteenable),  //                                             .byteenable
		.nios2_gen2_0_debug_mem_slave_waitrequest           (mm_interconnect_0_nios2_gen2_0_debug_mem_slave_waitrequest), //                                             .waitrequest
		.nios2_gen2_0_debug_mem_slave_debugaccess           (mm_interconnect_0_nios2_gen2_0_debug_mem_slave_debugaccess), //                                             .debugaccess
		.onchip_memory2_s1_address                          (mm_interconnect_0_onchip_memory2_s1_address),                //                            onchip_memory2_s1.address
		.onchip_memory2_s1_write                            (mm_interconnect_0_onchip_memory2_s1_write),                  //                                             .write
		.onchip_memory2_s1_readdata                         (mm_interconnect_0_onchip_memory2_s1_readdata),               //                                             .readdata
		.onchip_memory2_s1_writedata                        (mm_interconnect_0_onchip_memory2_s1_writedata),              //                                             .writedata
		.onchip_memory2_s1_byteenable                       (mm_interconnect_0_onchip_memory2_s1_byteenable),             //                                             .byteenable
		.onchip_memory2_s1_chipselect                       (mm_interconnect_0_onchip_memory2_s1_chipselect),             //                                             .chipselect
		.onchip_memory2_s1_clken                            (mm_interconnect_0_onchip_memory2_s1_clken),                  //                                             .clken
		.sdram_s1_address                                   (mm_interconnect_0_sdram_s1_address),                         //                                     sdram_s1.address
		.sdram_s1_write                                     (mm_interconnect_0_sdram_s1_write),                           //                                             .write
		.sdram_s1_read                                      (mm_interconnect_0_sdram_s1_read),                            //                                             .read
		.sdram_s1_readdata                                  (mm_interconnect_0_sdram_s1_readdata),                        //                                             .readdata
		.sdram_s1_writedata                                 (mm_interconnect_0_sdram_s1_writedata),                       //                                             .writedata
		.sdram_s1_byteenable                                (mm_interconnect_0_sdram_s1_byteenable),                      //                                             .byteenable
		.sdram_s1_readdatavalid                             (mm_interconnect_0_sdram_s1_readdatavalid),                   //                                             .readdatavalid
		.sdram_s1_waitrequest                               (mm_interconnect_0_sdram_s1_waitrequest),                     //                                             .waitrequest
		.sdram_s1_chipselect                                (mm_interconnect_0_sdram_s1_chipselect),                      //                                             .chipselect
		.sysid_qsys_control_slave_address                   (mm_interconnect_0_sysid_qsys_control_slave_address),         //                     sysid_qsys_control_slave.address
		.sysid_qsys_control_slave_readdata                  (mm_interconnect_0_sysid_qsys_control_slave_readdata),        //                                             .readdata
		.timer_s1_address                                   (mm_interconnect_0_timer_s1_address),                         //                                     timer_s1.address
		.timer_s1_write                                     (mm_interconnect_0_timer_s1_write),                           //                                             .write
		.timer_s1_readdata                                  (mm_interconnect_0_timer_s1_readdata),                        //                                             .readdata
		.timer_s1_writedata                                 (mm_interconnect_0_timer_s1_writedata),                       //                                             .writedata
		.timer_s1_chipselect                                (mm_interconnect_0_timer_s1_chipselect)                       //                                             .chipselect
	);

	audio_nios_mm_interconnect_1 mm_interconnect_1 (
		.pll_outclk2_clk                                            (pll_outclk2_clk),                               //                                          pll_outclk2.clk
		.cpu_peripheral_bridge_m0_reset_reset_bridge_in_reset_reset (rst_controller_001_reset_out_reset),            // cpu_peripheral_bridge_m0_reset_reset_bridge_in_reset.reset
		.cpu_peripheral_bridge_m0_address                           (cpu_peripheral_bridge_m0_address),              //                             cpu_peripheral_bridge_m0.address
		.cpu_peripheral_bridge_m0_waitrequest                       (cpu_peripheral_bridge_m0_waitrequest),          //                                                     .waitrequest
		.cpu_peripheral_bridge_m0_burstcount                        (cpu_peripheral_bridge_m0_burstcount),           //                                                     .burstcount
		.cpu_peripheral_bridge_m0_byteenable                        (cpu_peripheral_bridge_m0_byteenable),           //                                                     .byteenable
		.cpu_peripheral_bridge_m0_read                              (cpu_peripheral_bridge_m0_read),                 //                                                     .read
		.cpu_peripheral_bridge_m0_readdata                          (cpu_peripheral_bridge_m0_readdata),             //                                                     .readdata
		.cpu_peripheral_bridge_m0_readdatavalid                     (cpu_peripheral_bridge_m0_readdatavalid),        //                                                     .readdatavalid
		.cpu_peripheral_bridge_m0_write                             (cpu_peripheral_bridge_m0_write),                //                                                     .write
		.cpu_peripheral_bridge_m0_writedata                         (cpu_peripheral_bridge_m0_writedata),            //                                                     .writedata
		.cpu_peripheral_bridge_m0_debugaccess                       (cpu_peripheral_bridge_m0_debugaccess),          //                                                     .debugaccess
		.i2c_scl_s1_address                                         (mm_interconnect_1_i2c_scl_s1_address),          //                                           i2c_scl_s1.address
		.i2c_scl_s1_write                                           (mm_interconnect_1_i2c_scl_s1_write),            //                                                     .write
		.i2c_scl_s1_readdata                                        (mm_interconnect_1_i2c_scl_s1_readdata),         //                                                     .readdata
		.i2c_scl_s1_writedata                                       (mm_interconnect_1_i2c_scl_s1_writedata),        //                                                     .writedata
		.i2c_scl_s1_chipselect                                      (mm_interconnect_1_i2c_scl_s1_chipselect),       //                                                     .chipselect
		.i2c_sda_s1_address                                         (mm_interconnect_1_i2c_sda_s1_address),          //                                           i2c_sda_s1.address
		.i2c_sda_s1_write                                           (mm_interconnect_1_i2c_sda_s1_write),            //                                                     .write
		.i2c_sda_s1_readdata                                        (mm_interconnect_1_i2c_sda_s1_readdata),         //                                                     .readdata
		.i2c_sda_s1_writedata                                       (mm_interconnect_1_i2c_sda_s1_writedata),        //                                                     .writedata
		.i2c_sda_s1_chipselect                                      (mm_interconnect_1_i2c_sda_s1_chipselect),       //                                                     .chipselect
		.key_s1_address                                             (mm_interconnect_1_key_s1_address),              //                                               key_s1.address
		.key_s1_write                                               (mm_interconnect_1_key_s1_write),                //                                                     .write
		.key_s1_readdata                                            (mm_interconnect_1_key_s1_readdata),             //                                                     .readdata
		.key_s1_writedata                                           (mm_interconnect_1_key_s1_writedata),            //                                                     .writedata
		.key_s1_chipselect                                          (mm_interconnect_1_key_s1_chipselect),           //                                                     .chipselect
		.pio_led_s1_address                                         (mm_interconnect_1_pio_led_s1_address),          //                                           pio_led_s1.address
		.pio_led_s1_write                                           (mm_interconnect_1_pio_led_s1_write),            //                                                     .write
		.pio_led_s1_readdata                                        (mm_interconnect_1_pio_led_s1_readdata),         //                                                     .readdata
		.pio_led_s1_writedata                                       (mm_interconnect_1_pio_led_s1_writedata),        //                                                     .writedata
		.pio_led_s1_chipselect                                      (mm_interconnect_1_pio_led_s1_chipselect),       //                                                     .chipselect
		.seg7_avalon_slave_address                                  (mm_interconnect_1_seg7_avalon_slave_address),   //                                    seg7_avalon_slave.address
		.seg7_avalon_slave_write                                    (mm_interconnect_1_seg7_avalon_slave_write),     //                                                     .write
		.seg7_avalon_slave_read                                     (mm_interconnect_1_seg7_avalon_slave_read),      //                                                     .read
		.seg7_avalon_slave_readdata                                 (mm_interconnect_1_seg7_avalon_slave_readdata),  //                                                     .readdata
		.seg7_avalon_slave_writedata                                (mm_interconnect_1_seg7_avalon_slave_writedata), //                                                     .writedata
		.sw_s1_address                                              (mm_interconnect_1_sw_s1_address),               //                                                sw_s1.address
		.sw_s1_write                                                (mm_interconnect_1_sw_s1_write),                 //                                                     .write
		.sw_s1_readdata                                             (mm_interconnect_1_sw_s1_readdata),              //                                                     .readdata
		.sw_s1_writedata                                            (mm_interconnect_1_sw_s1_writedata),             //                                                     .writedata
		.sw_s1_chipselect                                           (mm_interconnect_1_sw_s1_chipselect)             //                                                     .chipselect
	);

	audio_nios_irq_mapper irq_mapper (
		.clk           (pll_outclk0_clk),                    //       clk.clk
		.reset         (rst_controller_003_reset_out_reset), // clk_reset.reset
		.receiver0_irq (irq_mapper_receiver0_irq),           // receiver0.irq
		.receiver1_irq (irq_mapper_receiver1_irq),           // receiver1.irq
		.receiver2_irq (irq_mapper_receiver2_irq),           // receiver2.irq
		.receiver3_irq (irq_mapper_receiver3_irq),           // receiver3.irq
		.sender_irq    (nios2_gen2_0_irq_irq)                //    sender.irq
	);

	altera_irq_clock_crosser #(
		.IRQ_WIDTH (1)
	) irq_synchronizer (
		.receiver_clk   (pll_outclk2_clk),                    //       receiver_clk.clk
		.sender_clk     (pll_outclk0_clk),                    //         sender_clk.clk
		.receiver_reset (rst_controller_001_reset_out_reset), // receiver_clk_reset.reset
		.sender_reset   (rst_controller_003_reset_out_reset), //   sender_clk_reset.reset
		.receiver_irq   (irq_synchronizer_receiver_irq),      //           receiver.irq
		.sender_irq     (irq_mapper_receiver2_irq)            //             sender.irq
	);

	altera_irq_clock_crosser #(
		.IRQ_WIDTH (1)
	) irq_synchronizer_001 (
		.receiver_clk   (pll_outclk2_clk),                    //       receiver_clk.clk
		.sender_clk     (pll_outclk0_clk),                    //         sender_clk.clk
		.receiver_reset (rst_controller_001_reset_out_reset), // receiver_clk_reset.reset
		.sender_reset   (rst_controller_003_reset_out_reset), //   sender_clk_reset.reset
		.receiver_irq   (irq_synchronizer_001_receiver_irq),  //           receiver.irq
		.sender_irq     (irq_mapper_receiver3_irq)            //             sender.irq
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (1),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (0),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller (
		.reset_in0      (~reset_reset_n),                 // reset_in0.reset
		.clk            (altpll_audio_outclk0_clk),       //       clk.clk
		.reset_out      (rst_controller_reset_out_reset), // reset_out.reset
		.reset_req      (),                               // (terminated)
		.reset_req_in0  (1'b0),                           // (terminated)
		.reset_in1      (1'b0),                           // (terminated)
		.reset_req_in1  (1'b0),                           // (terminated)
		.reset_in2      (1'b0),                           // (terminated)
		.reset_req_in2  (1'b0),                           // (terminated)
		.reset_in3      (1'b0),                           // (terminated)
		.reset_req_in3  (1'b0),                           // (terminated)
		.reset_in4      (1'b0),                           // (terminated)
		.reset_req_in4  (1'b0),                           // (terminated)
		.reset_in5      (1'b0),                           // (terminated)
		.reset_req_in5  (1'b0),                           // (terminated)
		.reset_in6      (1'b0),                           // (terminated)
		.reset_req_in6  (1'b0),                           // (terminated)
		.reset_in7      (1'b0),                           // (terminated)
		.reset_req_in7  (1'b0),                           // (terminated)
		.reset_in8      (1'b0),                           // (terminated)
		.reset_req_in8  (1'b0),                           // (terminated)
		.reset_in9      (1'b0),                           // (terminated)
		.reset_req_in9  (1'b0),                           // (terminated)
		.reset_in10     (1'b0),                           // (terminated)
		.reset_req_in10 (1'b0),                           // (terminated)
		.reset_in11     (1'b0),                           // (terminated)
		.reset_req_in11 (1'b0),                           // (terminated)
		.reset_in12     (1'b0),                           // (terminated)
		.reset_req_in12 (1'b0),                           // (terminated)
		.reset_in13     (1'b0),                           // (terminated)
		.reset_req_in13 (1'b0),                           // (terminated)
		.reset_in14     (1'b0),                           // (terminated)
		.reset_req_in14 (1'b0),                           // (terminated)
		.reset_in15     (1'b0),                           // (terminated)
		.reset_req_in15 (1'b0)                            // (terminated)
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (1),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (0),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller_001 (
		.reset_in0      (~reset_reset_n),                     // reset_in0.reset
		.clk            (pll_outclk2_clk),                    //       clk.clk
		.reset_out      (rst_controller_001_reset_out_reset), // reset_out.reset
		.reset_req      (),                                   // (terminated)
		.reset_req_in0  (1'b0),                               // (terminated)
		.reset_in1      (1'b0),                               // (terminated)
		.reset_req_in1  (1'b0),                               // (terminated)
		.reset_in2      (1'b0),                               // (terminated)
		.reset_req_in2  (1'b0),                               // (terminated)
		.reset_in3      (1'b0),                               // (terminated)
		.reset_req_in3  (1'b0),                               // (terminated)
		.reset_in4      (1'b0),                               // (terminated)
		.reset_req_in4  (1'b0),                               // (terminated)
		.reset_in5      (1'b0),                               // (terminated)
		.reset_req_in5  (1'b0),                               // (terminated)
		.reset_in6      (1'b0),                               // (terminated)
		.reset_req_in6  (1'b0),                               // (terminated)
		.reset_in7      (1'b0),                               // (terminated)
		.reset_req_in7  (1'b0),                               // (terminated)
		.reset_in8      (1'b0),                               // (terminated)
		.reset_req_in8  (1'b0),                               // (terminated)
		.reset_in9      (1'b0),                               // (terminated)
		.reset_req_in9  (1'b0),                               // (terminated)
		.reset_in10     (1'b0),                               // (terminated)
		.reset_req_in10 (1'b0),                               // (terminated)
		.reset_in11     (1'b0),                               // (terminated)
		.reset_req_in11 (1'b0),                               // (terminated)
		.reset_in12     (1'b0),                               // (terminated)
		.reset_req_in12 (1'b0),                               // (terminated)
		.reset_in13     (1'b0),                               // (terminated)
		.reset_req_in13 (1'b0),                               // (terminated)
		.reset_in14     (1'b0),                               // (terminated)
		.reset_req_in14 (1'b0),                               // (terminated)
		.reset_in15     (1'b0),                               // (terminated)
		.reset_req_in15 (1'b0)                                // (terminated)
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (1),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (1),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller_002 (
		.reset_in0      (~reset_reset_n),                         // reset_in0.reset
		.clk            (pll_outclk0_clk),                        //       clk.clk
		.reset_out      (rst_controller_002_reset_out_reset),     // reset_out.reset
		.reset_req      (rst_controller_002_reset_out_reset_req), //          .reset_req
		.reset_req_in0  (1'b0),                                   // (terminated)
		.reset_in1      (1'b0),                                   // (terminated)
		.reset_req_in1  (1'b0),                                   // (terminated)
		.reset_in2      (1'b0),                                   // (terminated)
		.reset_req_in2  (1'b0),                                   // (terminated)
		.reset_in3      (1'b0),                                   // (terminated)
		.reset_req_in3  (1'b0),                                   // (terminated)
		.reset_in4      (1'b0),                                   // (terminated)
		.reset_req_in4  (1'b0),                                   // (terminated)
		.reset_in5      (1'b0),                                   // (terminated)
		.reset_req_in5  (1'b0),                                   // (terminated)
		.reset_in6      (1'b0),                                   // (terminated)
		.reset_req_in6  (1'b0),                                   // (terminated)
		.reset_in7      (1'b0),                                   // (terminated)
		.reset_req_in7  (1'b0),                                   // (terminated)
		.reset_in8      (1'b0),                                   // (terminated)
		.reset_req_in8  (1'b0),                                   // (terminated)
		.reset_in9      (1'b0),                                   // (terminated)
		.reset_req_in9  (1'b0),                                   // (terminated)
		.reset_in10     (1'b0),                                   // (terminated)
		.reset_req_in10 (1'b0),                                   // (terminated)
		.reset_in11     (1'b0),                                   // (terminated)
		.reset_req_in11 (1'b0),                                   // (terminated)
		.reset_in12     (1'b0),                                   // (terminated)
		.reset_req_in12 (1'b0),                                   // (terminated)
		.reset_in13     (1'b0),                                   // (terminated)
		.reset_req_in13 (1'b0),                                   // (terminated)
		.reset_in14     (1'b0),                                   // (terminated)
		.reset_req_in14 (1'b0),                                   // (terminated)
		.reset_in15     (1'b0),                                   // (terminated)
		.reset_req_in15 (1'b0)                                    // (terminated)
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (2),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (1),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller_003 (
		.reset_in0      (~reset_reset_n),                         // reset_in0.reset
		.reset_in1      (nios2_gen2_0_debug_reset_request_reset), // reset_in1.reset
		.clk            (pll_outclk0_clk),                        //       clk.clk
		.reset_out      (rst_controller_003_reset_out_reset),     // reset_out.reset
		.reset_req      (rst_controller_003_reset_out_reset_req), //          .reset_req
		.reset_req_in0  (1'b0),                                   // (terminated)
		.reset_req_in1  (1'b0),                                   // (terminated)
		.reset_in2      (1'b0),                                   // (terminated)
		.reset_req_in2  (1'b0),                                   // (terminated)
		.reset_in3      (1'b0),                                   // (terminated)
		.reset_req_in3  (1'b0),                                   // (terminated)
		.reset_in4      (1'b0),                                   // (terminated)
		.reset_req_in4  (1'b0),                                   // (terminated)
		.reset_in5      (1'b0),                                   // (terminated)
		.reset_req_in5  (1'b0),                                   // (terminated)
		.reset_in6      (1'b0),                                   // (terminated)
		.reset_req_in6  (1'b0),                                   // (terminated)
		.reset_in7      (1'b0),                                   // (terminated)
		.reset_req_in7  (1'b0),                                   // (terminated)
		.reset_in8      (1'b0),                                   // (terminated)
		.reset_req_in8  (1'b0),                                   // (terminated)
		.reset_in9      (1'b0),                                   // (terminated)
		.reset_req_in9  (1'b0),                                   // (terminated)
		.reset_in10     (1'b0),                                   // (terminated)
		.reset_req_in10 (1'b0),                                   // (terminated)
		.reset_in11     (1'b0),                                   // (terminated)
		.reset_req_in11 (1'b0),                                   // (terminated)
		.reset_in12     (1'b0),                                   // (terminated)
		.reset_req_in12 (1'b0),                                   // (terminated)
		.reset_in13     (1'b0),                                   // (terminated)
		.reset_req_in13 (1'b0),                                   // (terminated)
		.reset_in14     (1'b0),                                   // (terminated)
		.reset_req_in14 (1'b0),                                   // (terminated)
		.reset_in15     (1'b0),                                   // (terminated)
		.reset_req_in15 (1'b0)                                    // (terminated)
	);

endmodule
